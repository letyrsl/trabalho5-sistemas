`include "bo.v"

module quadratic_eq(
  input[7:0] x,
  input[15:0] a,
  input[15:0] b,
  input[15:0] c,
  input inicio,
  input clock,
  input reset,

  output pronto,
  output[15:0] resultado
);
  // bo bo_0(x, a, b, c, );
endmodule